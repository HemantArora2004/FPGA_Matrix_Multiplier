`timescale 1ns / 1ps
module Matrix_Multiplier(

    );
endmodule
