`timescale 1ns / 1ps
module axi_stream_slave(
    input logic clk,
    input logic reset,
    input logic s_axis_valid,
    output logic s_axis_ready,
    input logic s_axis_data,
    input logic s_axis_last
);


endmodule
